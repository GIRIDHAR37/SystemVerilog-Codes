class example;
  
  rand bit [7:0]a[3][3][3];
  
  constraint a_c{
    foreach(a[i,j,k]){
      foreach(a[x,y,z]){
        if((i!=x)||(j!=y)||(k!=z))
          a[i][j][k]!=a[x][y][z];
      }
    }
  }
  
  function void print();
    $display("Array a elements : %p",a);
  endfunction
  
endclass

module top;
  
  example ex=new();
  
  initial begin
    repeat(10) begin
      ex.randomize();
      ex.print();
    end
  end
  
endmodule

// output :

/*
# Array a elements : '{'{'{213, 159, 188}, '{168, 147, 236}, '{203, 24, 7}}, '{'{73, 193, 224}, '{205, 91, 180}, '{37, 173, 52}}, '{'{26, 148, 190}, '{11, 166, 45}, '{136, 54, 158}}}
# Array a elements : '{'{'{31, 58, 153}, '{120, 211, 179}, '{40, 47, 93}}, '{'{63, 224, 51}, '{123, 52, 57}, '{187, 175, 142}}, '{'{68, 79, 65}, '{36, 133, 131}, '{176, 111, 49}}}
# Array a elements : '{'{'{164, 204, 25}, '{23, 173, 230}, '{152, 56, 213}}, '{'{79, 82, 148}, '{212, 196, 21}, '{143, 116, 77}}, '{'{72, 86, 169}, '{34, 226, 180}, '{62, 174, 39}}}
# Array a elements : '{'{'{223, 162, 225}, '{62, 255, 24}, '{164, 153, 27}}, '{'{159, 126, 227}, '{41, 47, 15}, '{75, 37, 178}}, '{'{35, 16, 7}, '{113, 222, 114}, '{34, 169, 84}}}
# Array a elements : '{'{'{199, 88, 235}, '{6, 101, 67}, '{103, 53, 193}}, '{'{181, 90, 207}, '{114, 213, 131}, '{157, 120, 36}}, '{'{24, 178, 19}, '{169, 248, 134}, '{58, 93, 23}}}
# Array a elements : '{'{'{54, 69, 41}, '{157, 21, 97}, '{249, 48, 131}}, '{'{226, 178, 242}, '{83, 100, 38}, '{2, 87, 188}}, '{'{151, 47, 170}, '{114, 183, 229}, '{46, 175, 174}}}
# Array a elements : '{'{'{15, 254, 23}, '{132, 101, 203}, '{113, 91, 169}}, '{'{200, 150, 249}, '{146, 166, 204}, '{148, 112, 96}}, '{'{185, 40, 245}, '{226, 54, 208}, '{238, 164, 56}}}
# Array a elements : '{'{'{5, 54, 98}, '{199, 91, 185}, '{192, 241, 187}}, '{'{219, 254, 62}, '{197, 73, 148}, '{141, 209, 247}}, '{'{243, 228, 111}, '{29, 64, 147}, '{181, 66, 252}}}
# Array a elements : '{'{'{111, 203, 108}, '{125, 134, 72}, '{201, 129, 25}}, '{'{46, 188, 205}, '{207, 64, 211}, '{172, 221, 194}}, '{'{114, 234, 21}, '{213, 216, 177}, '{33, 49, 118}}}
# Array a elements : '{'{'{87, 114, 202}, '{218, 221, 251}, '{204, 217, 27}}, '{'{158, 177, 167}, '{124, 76, 215}, '{46, 102, 143}}, '{'{12, 222, 39}, '{136, 110, 226}, '{106, 228, 234}}}
*/

